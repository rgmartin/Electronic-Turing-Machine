CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 0 22 70 10
176 79 1598 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
42991632 0
0
6 Title:
5 Name:
0
0
0
196
13 Logic Switch~
5 292 114 0 1 11
0 41
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
41410.4 0
0
13 Logic Switch~
5 316 114 0 1 11
0 40
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
41410.4 1
0
13 Logic Switch~
5 340 113 0 1 11
0 39
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
41410.4 2
0
13 Logic Switch~
5 363 111 0 1 11
0 38
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
41410.4 3
0
13 Logic Switch~
5 386 112 0 1 11
0 37
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
41410.4 4
0
13 Logic Switch~
5 431 112 0 1 11
0 35
0
0 0 20592 270
2 0V
-7 -22 7 -14
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
41410.4 5
0
13 Logic Switch~
5 453 112 0 1 11
0 34
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
41410.4 6
0
13 Logic Switch~
5 476 112 0 1 11
0 33
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
41410.4 7
0
13 Logic Switch~
5 498 111 0 1 11
0 32
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
41410.4 8
0
13 Logic Switch~
5 520 111 0 1 11
0 31
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
41410.4 9
0
13 Logic Switch~
5 543 109 0 1 11
0 30
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
41410.4 10
0
13 Logic Switch~
5 566 110 0 1 11
0 29
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
41410.4 11
0
13 Logic Switch~
5 591 109 0 1 11
0 28
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
41410.4 12
0
13 Logic Switch~
5 614 111 0 1 11
0 27
0
0 0 20592 270
2 0V
-6 -21 8 -13
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
41410.4 13
0
13 Logic Switch~
5 638 111 0 1 11
0 26
0
0 0 20592 270
2 0V
-6 -21 8 -13
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
41410.4 14
0
13 Logic Switch~
5 410 113 0 1 11
0 36
0
0 0 20720 270
2 0V
-7 -22 7 -14
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
41410.4 15
0
13 Logic Switch~
5 348 397 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-7 -22 7 -14
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5616 0 0
2
41410.4 16
0
13 Logic Switch~
5 283 397 0 1 11
0 46
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
41410.4 17
0
13 Logic Switch~
5 305 398 0 1 11
0 45
0
0 0 20592 270
2 0V
-7 -22 7 -14
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
41410.4 18
0
13 Logic Switch~
5 327 396 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-7 -22 7 -14
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3108 0 0
2
41410.4 19
0
13 Logic Switch~
5 234 664 0 1 11
0 42
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4299 0 0
2
41410.4 20
0
9 Inverter~
13 1074 860 0 2 22
0 42 4
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U68B
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 44 0
1 U
9672 0 0
2
41410.4 21
0
9 Inverter~
13 268 565 0 2 22
0 42 25
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U68A
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 44 0
1 U
7876 0 0
2
41410.4 22
0
10 Buffer 3S~
219 293 136 0 3 22
0 41 25 24
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U63A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 39 0
1 U
6369 0 0
2
41410.4 23
0
10 Buffer 3S~
219 317 136 0 3 22
0 40 25 23
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U63B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 39 0
1 U
9172 0 0
2
41410.4 24
0
10 Buffer 3S~
219 341 135 0 3 22
0 39 25 22
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U63C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 39 0
1 U
7100 0 0
2
41410.4 25
0
10 Buffer 3S~
219 365 134 0 3 22
0 38 25 21
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U63D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 39 0
1 U
3820 0 0
2
41410.4 26
0
10 Buffer 3S~
219 387 134 0 3 22
0 37 25 20
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U64A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 40 0
1 U
7678 0 0
2
41410.4 27
0
10 Buffer 3S~
219 410 134 0 3 22
0 36 25 19
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U64B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 40 0
1 U
961 0 0
2
41410.4 28
0
10 Buffer 3S~
219 432 135 0 3 22
0 35 25 18
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U64C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 40 0
1 U
3178 0 0
2
41410.4 29
0
10 Buffer 3S~
219 454 135 0 3 22
0 34 25 17
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U64D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 40 0
1 U
3409 0 0
2
41410.4 30
0
10 Buffer 3S~
219 478 135 0 3 22
0 33 25 16
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U65A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
3951 0 0
2
41410.4 31
0
10 Buffer 3S~
219 500 134 0 3 22
0 32 25 15
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U65B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 41 0
1 U
8885 0 0
2
41410.4 32
0
10 Buffer 3S~
219 521 134 0 3 22
0 31 25 14
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U65C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 41 0
1 U
3780 0 0
2
41410.4 33
0
10 Buffer 3S~
219 544 135 0 3 22
0 30 25 13
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U65D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 41 0
1 U
9265 0 0
2
41410.4 34
0
10 Buffer 3S~
219 567 135 0 3 22
0 29 25 12
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U66A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 42 0
1 U
9442 0 0
2
41410.4 35
0
10 Buffer 3S~
219 592 135 0 3 22
0 28 25 11
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U66B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 42 0
1 U
9424 0 0
2
41410.4 36
0
10 Buffer 3S~
219 615 135 0 3 22
0 27 25 10
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U66C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 42 0
1 U
9968 0 0
2
41410.4 37
0
10 Buffer 3S~
219 639 135 0 3 22
0 26 25 9
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U66D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 42 0
1 U
9281 0 0
2
41410.4 38
0
10 Buffer 3S~
219 348 421 0 3 22
0 43 25 7
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U67D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 43 0
1 U
8464 0 0
2
41410.4 39
0
10 Buffer 3S~
219 327 421 0 3 22
0 44 25 6
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U67C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 43 0
1 U
7168 0 0
2
41410.4 40
0
10 Buffer 3S~
219 306 421 0 3 22
0 45 25 5
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U67B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 43 0
1 U
3171 0 0
2
41410.4 41
0
10 Buffer 3S~
219 285 421 0 3 22
0 46 25 8
0
0 0 112 782
8 BUFFER3S
-27 -51 29 -43
4 U67A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 43 0
1 U
4139 0 0
2
41410.4 42
0
7 Ground~
168 787 715 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
41410.4 43
0
11 SUM-REST-4B
94 2023 747 0 10 21
0 114 113 112 111 122 123 108 121 110
107
11 SUM-REST-4B
1 0 4240 0
0
3 U39
-5 -62 16 -54
0
0
0
0
0
0
21

0 1 2 3 4 5 6 9 10 11
12 1 2 3 4 5 6 9 10 11
12 0
0 0 0 0 1 0 0 0
1 U
5283 0 0
2
5.89615e-315 0
0
9 Inverter~
13 989 225 0 2 22
0 23 153
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U1D
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6874 0 0
2
5.89615e-315 5.26354e-315
0
14 Logic Display~
6 974 148 0 1 2
10 101
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L2
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.89615e-315 5.30499e-315
0
13 SR Flip-Flop~
219 980 212 0 4 9
0 23 153 212 101
0
0 0 4464 90
4 0001
-11 -29 17 -21
2 U3
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.89615e-315 5.32571e-315
0
9 Inverter~
13 886 228 0 2 22
0 24 154
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U1C
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
969 0 0
2
5.89615e-315 5.34643e-315
0
14 Logic Display~
6 871 151 0 1 2
10 102
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89615e-315 5.3568e-315
0
13 SR Flip-Flop~
219 877 215 0 4 9
0 24 154 213 102
0
0 0 4464 90
4 0000
-11 -29 17 -21
2 U2
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3751 0 0
2
5.89615e-315 5.36716e-315
0
9 Inverter~
13 1094 226 0 2 22
0 22 155
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U1E
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
4292 0 0
2
5.89615e-315 5.37752e-315
0
14 Logic Display~
6 1079 149 0 1 2
10 100
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89615e-315 5.38788e-315
0
13 SR Flip-Flop~
219 1085 213 0 4 9
0 22 155 214 100
0
0 0 4464 90
4 0010
-11 -29 17 -21
2 U4
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.89615e-315 5.39306e-315
0
13 SR Flip-Flop~
219 1200 212 0 4 9
0 21 156 215 98
0
0 0 4464 90
4 0011
-11 -29 17 -21
2 U8
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6357 0 0
2
5.89615e-315 5.39824e-315
0
14 Logic Display~
6 1194 148 0 1 2
10 98
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L6
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
5.89615e-315 5.40342e-315
0
9 Inverter~
13 1209 225 0 2 22
0 21 156
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7B
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3976 0 0
2
5.89615e-315 5.4086e-315
0
9 Inverter~
13 1313 223 0 2 22
0 20 157
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7A
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7634 0 0
2
5.89615e-315 5.41378e-315
0
14 Logic Display~
6 1298 146 0 1 2
10 99
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L5
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.89615e-315 5.41896e-315
0
13 SR Flip-Flop~
219 1304 210 0 4 9
0 20 157 216 99
0
0 0 4464 90
4 0100
-11 -29 17 -21
2 U6
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6748 0 0
2
5.89615e-315 5.42414e-315
0
13 SR Flip-Flop~
219 1412 210 0 4 9
0 19 158 217 97
0
0 0 4464 90
4 0101
-11 -29 17 -21
2 U5
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6901 0 0
2
5.89615e-315 5.42933e-315
0
14 Logic Display~
6 1406 146 0 1 2
10 97
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L4
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
5.89615e-315 5.43192e-315
0
9 Inverter~
13 1421 223 0 2 22
0 19 158
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U1F
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3277 0 0
2
5.89615e-315 5.43451e-315
0
9 Inverter~
13 1530 223 0 2 22
0 18 159
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U14B
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
4212 0 0
2
5.89615e-315 5.4371e-315
0
14 Logic Display~
6 1515 146 0 1 2
10 96
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L12
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.89615e-315 5.43969e-315
0
13 SR Flip-Flop~
219 1521 210 0 4 9
0 18 159 218 96
0
0 0 4464 90
4 0110
-11 -29 17 -21
3 U15
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5551 0 0
2
5.89615e-315 5.44228e-315
0
13 SR Flip-Flop~
219 1629 211 0 4 9
0 17 161 219 95
0
0 0 4464 90
4 0111
-11 -29 17 -21
3 U13
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
5.89615e-315 5.44487e-315
0
14 Logic Display~
6 1623 147 0 1 2
10 95
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L11
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.89615e-315 5.44746e-315
0
9 Inverter~
13 1638 224 0 2 22
0 17 161
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U14A
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9592 0 0
2
5.89615e-315 5.45005e-315
0
13 SR Flip-Flop~
219 1732 211 0 4 9
0 16 160 220 94
0
0 0 4464 90
4 1000
-11 -29 17 -21
3 U12
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8748 0 0
2
5.89615e-315 5.45264e-315
0
14 Logic Display~
6 1726 147 0 1 2
10 94
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L10
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89615e-315 5.45523e-315
0
9 Inverter~
13 1741 224 0 2 22
0 16 160
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7F
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
631 0 0
2
5.89615e-315 5.45782e-315
0
9 Inverter~
13 1851 222 0 2 22
0 15 152
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7C
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9466 0 0
2
5.89615e-315 5.46041e-315
0
14 Logic Display~
6 1836 145 0 1 2
10 93
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L7
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
5.89615e-315 5.463e-315
0
13 SR Flip-Flop~
219 1842 209 0 4 9
0 15 152 221 93
0
0 0 4464 90
4 1001
-11 -29 17 -21
2 U9
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7693 0 0
2
5.89615e-315 5.46559e-315
0
13 SR Flip-Flop~
219 1948 212 0 4 9
0 14 146 222 92
0
0 0 4464 90
4 1010
-11 -29 17 -21
3 U10
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3723 0 0
2
5.89615e-315 5.46818e-315
0
14 Logic Display~
6 1942 148 0 1 2
10 92
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L8
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.89615e-315 5.47077e-315
0
9 Inverter~
13 1957 225 0 2 22
0 14 146
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7D
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
6263 0 0
2
5.89615e-315 0
0
9 Inverter~
13 2064 224 0 2 22
0 13 147
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U7E
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
4900 0 0
2
5.89615e-315 5.26354e-315
0
14 Logic Display~
6 2049 147 0 1 2
10 91
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L9
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
5.89615e-315 5.30499e-315
0
13 SR Flip-Flop~
219 2055 211 0 4 9
0 13 147 223 91
0
0 0 4464 90
4 1011
-11 -29 17 -21
3 U11
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3221 0 0
2
5.89615e-315 5.32571e-315
0
13 SR Flip-Flop~
219 2169 212 0 4 9
0 12 148 224 90
0
0 0 4464 90
4 1100
-11 -29 17 -21
3 U20
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3215 0 0
2
5.89615e-315 5.34643e-315
0
14 Logic Display~
6 2163 148 0 1 2
10 90
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L17
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
5.89615e-315 5.3568e-315
0
9 Inverter~
13 2178 225 0 2 22
0 12 148
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U21A
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7121 0 0
2
5.89615e-315 5.36716e-315
0
9 Inverter~
13 2299 223 0 2 22
0 11 149
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U14F
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
4484 0 0
2
5.89615e-315 5.37752e-315
0
14 Logic Display~
6 2284 146 0 1 2
10 89
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L16
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.89615e-315 5.38788e-315
0
13 SR Flip-Flop~
219 2290 210 0 4 9
0 11 149 225 89
0
0 0 4464 90
4 1101
-11 -29 17 -21
3 U19
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7804 0 0
2
5.89615e-315 5.39306e-315
0
13 SR Flip-Flop~
219 2402 210 0 4 9
0 10 150 226 88
0
0 0 4464 90
4 1110
-11 -29 17 -21
3 U16
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5523 0 0
2
5.89615e-315 5.39824e-315
0
14 Logic Display~
6 2396 146 0 1 2
10 88
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L13
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.89615e-315 5.40342e-315
0
9 Inverter~
13 2411 223 0 2 22
0 10 150
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U14C
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3465 0 0
2
5.89615e-315 5.4086e-315
0
13 SR Flip-Flop~
219 2523 208 0 4 9
0 9 151 227 87
0
0 0 4464 90
4 1111
-11 -29 17 -21
3 U17
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8396 0 0
2
5.89615e-315 5.41378e-315
0
14 Logic Display~
6 2517 144 0 1 2
10 87
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 L14
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.89615e-315 5.41896e-315
0
9 Inverter~
13 2532 221 0 2 22
0 9 151
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U14D
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
7849 0 0
2
5.89615e-315 5.42414e-315
0
10 Buffer 3S~
219 871 267 0 3 22
0 67 145 24
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U33A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6343 0 0
2
5.89615e-315 5.42933e-315
0
10 Buffer 3S~
219 974 262 0 3 22
0 67 143 23
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U33B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7376 0 0
2
5.89615e-315 5.43192e-315
0
10 Buffer 3S~
219 1079 262 0 3 22
0 67 142 22
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U33C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
9156 0 0
2
5.89615e-315 5.43451e-315
0
10 Buffer 3S~
219 1194 262 0 3 22
0 67 144 21
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U33D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
5776 0 0
2
5.89615e-315 5.4371e-315
0
10 Buffer 3S~
219 1298 262 0 3 22
0 67 141 20
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U25A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7207 0 0
2
5.89615e-315 5.43969e-315
0
10 Buffer 3S~
219 1406 260 0 3 22
0 67 140 19
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U26A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4459 0 0
2
5.89615e-315 5.44228e-315
0
10 Buffer 3S~
219 1515 261 0 3 22
0 67 139 18
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U27A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3760 0 0
2
5.89615e-315 5.44487e-315
0
10 Buffer 3S~
219 1623 261 0 3 22
0 67 115 17
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U28A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
754 0 0
2
5.89615e-315 5.44746e-315
0
10 Buffer 3S~
219 1726 265 0 3 22
0 67 138 16
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U34A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
9767 0 0
2
5.89615e-315 5.45005e-315
0
10 Buffer 3S~
219 1836 261 0 3 22
0 67 137 15
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U34B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
7978 0 0
2
5.89615e-315 5.45264e-315
0
10 Buffer 3S~
219 1942 264 0 3 22
0 67 136 14
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U34C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
3142 0 0
2
5.89615e-315 5.45523e-315
0
10 Buffer 3S~
219 2164 263 0 3 22
0 67 134 12
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U35A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
3284 0 0
2
5.89615e-315 5.45782e-315
0
10 Buffer 3S~
219 2284 261 0 3 22
0 67 133 11
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U35B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
659 0 0
2
5.89615e-315 5.46041e-315
0
10 Buffer 3S~
219 2396 263 0 3 22
0 67 132 10
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U35C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
3800 0 0
2
5.89615e-315 5.463e-315
0
10 Buffer 3S~
219 2517 262 0 3 22
0 67 131 9
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U35D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
6792 0 0
2
5.89615e-315 5.46559e-315
0
9 4-In AND~
219 901 457 0 5 22
0 70 126 125 124 84
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U36A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 16 0
1 U
3701 0 0
2
5.89615e-315 5.46818e-315
0
9 4-In AND~
219 1228 452 0 5 22
0 114 113 125 124 82
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U36B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 16 0
1 U
6316 0 0
2
5.89615e-315 5.47077e-315
0
9 4-In AND~
219 1006 456 0 5 22
0 114 126 125 124 83
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U37A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 17 0
1 U
8734 0 0
2
5.89615e-315 5.47207e-315
0
9 4-In AND~
219 1112 452 0 5 22
0 70 113 125 124 81
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U37B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 17 0
1 U
7988 0 0
2
5.89615e-315 5.47336e-315
0
9 4-In AND~
219 1441 450 0 5 22
0 114 126 112 124 78
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U38A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 18 0
1 U
3217 0 0
2
5.89615e-315 5.47466e-315
0
9 4-In AND~
219 1333 450 0 5 22
0 70 126 112 124 80
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U38B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 18 0
1 U
3965 0 0
2
5.89615e-315 5.47595e-315
0
9 4-In AND~
219 1551 447 0 5 22
0 70 113 112 124 79
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U40A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 20 0
1 U
8239 0 0
2
5.89615e-315 5.47725e-315
0
9 4-In AND~
219 2430 440 0 5 22
0 70 113 112 111 69
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U41A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 21 0
1 U
828 0 0
2
5.89615e-315 5.47854e-315
0
9 4-In AND~
219 1977 440 0 5 22
0 70 113 125 111 74
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U41B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 21 0
1 U
6187 0 0
2
5.89615e-315 5.47984e-315
0
9 4-In AND~
219 2084 438 0 5 22
0 114 113 125 111 73
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U42A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 22 0
1 U
7107 0 0
2
5.89615e-315 5.48113e-315
0
9 4-In AND~
219 1870 442 0 5 22
0 114 126 125 111 75
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U43A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 23 0
1 U
6433 0 0
2
5.89615e-315 5.48243e-315
0
9 4-In AND~
219 2198 442 0 5 22
0 70 126 112 111 72
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U43B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 23 0
1 U
8559 0 0
2
5.89615e-315 5.48372e-315
0
9 4-In AND~
219 1659 445 0 5 22
0 114 113 112 124 77
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U44A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 24 0
1 U
3674 0 0
2
5.89615e-315 5.48502e-315
0
9 4-In AND~
219 1762 450 0 5 22
0 70 126 125 111 76
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U44B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 24 0
1 U
5697 0 0
2
5.89615e-315 5.48631e-315
0
9 4-In AND~
219 2552 430 0 5 22
0 114 113 112 111 68
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U45A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 25 0
1 U
3805 0 0
2
5.89615e-315 5.48761e-315
0
9 4-In AND~
219 2318 435 0 5 22
0 114 126 112 111 71
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U45B
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 25 0
1 U
5219 0 0
2
5.89615e-315 5.4889e-315
0
13 SR Flip-Flop~
219 2658 589 0 4 9
0 7 130 70 114
0
0 0 4464 90
2 P1
-5 -26 9 -18
3 U18
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3795 0 0
2
5.89615e-315 5.4902e-315
0
9 Inverter~
13 2667 602 0 2 22
0 7 130
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U21B
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3637 0 0
2
5.89615e-315 5.49149e-315
0
9 Inverter~
13 2721 600 0 2 22
0 6 129
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U21C
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3226 0 0
2
5.89615e-315 5.49279e-315
0
13 SR Flip-Flop~
219 2712 587 0 4 9
0 6 129 126 113
0
0 0 4464 90
2 P2
-5 -29 9 -21
3 U22
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
6966 0 0
2
5.89615e-315 5.49408e-315
0
13 SR Flip-Flop~
219 2765 587 0 4 9
0 5 128 125 112
0
0 0 4464 90
2 P3
-4 -29 10 -21
3 U23
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9796 0 0
2
5.89615e-315 5.49538e-315
0
9 Inverter~
13 2774 600 0 2 22
0 5 128
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U21D
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
5952 0 0
2
5.89615e-315 5.49667e-315
0
9 Inverter~
13 2825 599 0 2 22
0 8 127
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U21E
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
3649 0 0
2
5.89615e-315 5.49797e-315
0
13 SR Flip-Flop~
219 2816 586 0 4 9
0 8 127 124 111
0
0 0 4464 90
2 P4
-4 -29 10 -21
3 U24
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3716 0 0
2
5.89615e-315 5.49926e-315
0
14 Logic Display~
6 1641 648 0 1 2
10 66
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 IB
-29 7 -15 15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
5.89615e-315 5.50056e-315
0
9 Inverter~
13 916 967 0 2 22
0 50 85
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4681 0 0
2
5.89615e-315 5.50185e-315
0
9 Inverter~
13 911 932 0 2 22
0 49 116
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9730 0 0
2
5.89615e-315 5.50315e-315
0
10 Buffer 3S~
219 1695 713 0 3 22
0 57 58 59
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U46A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
9874 0 0
2
5.89615e-315 5.50444e-315
0
10 Buffer 3S~
219 1695 771 0 3 22
0 56 58 122
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U46B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
364 0 0
2
5.89615e-315 5.50574e-315
0
10 Buffer 3S~
219 1695 822 0 3 22
0 55 58 123
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U46C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
3656 0 0
2
5.89615e-315 5.50703e-315
0
9 2-In AND~
219 1696 880 0 3 22
0 116 85 58
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U47A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 27 0
1 U
3131 0 0
2
5.89615e-315 5.50833e-315
0
13 SR Flip-Flop~
219 2301 685 0 4 9
0 103 65 228 120
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
3 NP1
-12 -32 9 -24
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6772 0 0
2
5.89615e-315 5.50963e-315
0
13 SR Flip-Flop~
219 2303 736 0 4 9
0 106 64 229 119
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
3 NP2
-10 -31 11 -23
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9557 0 0
2
5.89615e-315 5.51092e-315
0
13 SR Flip-Flop~
219 2305 791 0 4 9
0 105 63 230 118
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
3 NP3
-10 -30 11 -22
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5789 0 0
2
5.89615e-315 5.51222e-315
0
9 Inverter~
13 2259 718 0 2 22
0 106 64
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U48A
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 19 0
1 U
7328 0 0
2
5.89615e-315 5.51286e-315
0
9 Inverter~
13 2257 667 0 2 22
0 103 65
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U48B
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 19 0
1 U
4799 0 0
2
5.89615e-315 5.51351e-315
0
9 Inverter~
13 2261 773 0 2 22
0 105 63
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U48C
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 19 0
1 U
9196 0 0
2
5.89615e-315 5.51416e-315
0
9 Inverter~
13 2264 823 0 2 22
0 104 62
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U48D
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 19 0
1 U
3857 0 0
2
5.89615e-315 5.51481e-315
0
13 SR Flip-Flop~
219 2308 841 0 4 9
0 104 62 231 109
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
3 NP4
-10 -30 11 -22
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7125 0 0
2
5.89615e-315 5.51545e-315
0
13 SR Flip-Flop~
219 1749 668 0 4 9
0 59 60 232 67
0
0 0 4720 90
4 SRFF
-14 -53 14 -45
2 OB
-3 -28 11 -20
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3641 0 0
2
5.89615e-315 5.5161e-315
0
9 Inverter~
13 1758 683 0 2 22
0 59 60
0
0 0 112 90
6 74LS04
-21 -19 21 -11
4 U48E
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 19 0
1 U
9821 0 0
2
5.89615e-315 5.51675e-315
0
10 Buffer 3S~
219 2371 649 0 3 22
0 120 117 7
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U49A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
3187 0 0
2
5.89615e-315 5.5174e-315
0
10 Buffer 3S~
219 2371 700 0 3 22
0 119 117 6
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U49B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
762 0 0
2
5.89615e-315 5.51804e-315
0
10 Buffer 3S~
219 2371 755 0 3 22
0 118 117 5
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U49C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
39 0 0
2
5.89615e-315 5.51869e-315
0
10 Buffer 3S~
219 2373 805 0 3 22
0 109 117 8
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U49D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
9450 0 0
2
5.89615e-315 5.51934e-315
0
9 2-In AND~
219 2374 883 0 3 22
0 50 116 117
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U47C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
3236 0 0
2
5.89615e-315 5.51999e-315
0
10 Buffer 3S~
219 2173 701 0 3 22
0 110 58 106
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U30A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3321 0 0
2
5.89615e-315 5.52063e-315
0
10 Buffer 3S~
219 2173 649 0 3 22
0 107 58 103
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U29A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
8879 0 0
2
5.89615e-315 5.52128e-315
0
10 Buffer 3S~
219 2173 755 0 3 22
0 121 58 105
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U31A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
5433 0 0
2
5.89615e-315 5.52193e-315
0
10 Buffer 3S~
219 2173 805 0 3 22
0 108 58 104
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
4 U32A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3679 0 0
2
5.89615e-315 5.52258e-315
0
10 Buffer 3S~
219 912 269 0 3 22
0 102 84 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U50A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
9342 0 0
2
5.89615e-315 5.52322e-315
0
10 Buffer 3S~
219 1017 268 0 3 22
0 101 83 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U56A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 35 0
1 U
3623 0 0
2
5.89615e-315 5.52387e-315
0
10 Buffer 3S~
219 1123 270 0 3 22
0 100 81 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U56B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 35 0
1 U
3722 0 0
2
5.89615e-315 5.52452e-315
0
10 Buffer 3S~
219 1344 269 0 3 22
0 99 80 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U56C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 35 0
1 U
8993 0 0
2
5.89615e-315 5.52517e-315
0
10 Buffer 3S~
219 1239 269 0 3 22
0 98 82 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U56D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 35 0
1 U
3723 0 0
2
5.89615e-315 5.52581e-315
0
10 Buffer 3S~
219 1452 267 0 3 22
0 97 78 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U57A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 36 0
1 U
6244 0 0
2
5.89615e-315 5.52646e-315
0
10 Buffer 3S~
219 1562 267 0 3 22
0 96 79 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U57B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 36 0
1 U
6421 0 0
2
5.89615e-315 5.52711e-315
0
10 Buffer 3S~
219 1670 267 0 3 22
0 95 77 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U57C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 36 0
1 U
7743 0 0
2
5.89615e-315 5.52776e-315
0
10 Buffer 3S~
219 1773 270 0 3 22
0 94 76 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U57D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 36 0
1 U
9840 0 0
2
5.89615e-315 5.52841e-315
0
10 Buffer 3S~
219 1881 267 0 3 22
0 93 75 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U58A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 37 0
1 U
6910 0 0
2
5.89615e-315 5.52905e-315
0
10 Buffer 3S~
219 1988 271 0 3 22
0 92 74 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U58B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 37 0
1 U
449 0 0
2
5.89615e-315 5.5297e-315
0
10 Buffer 3S~
219 2095 270 0 3 22
0 91 73 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U58C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 37 0
1 U
8761 0 0
2
5.89615e-315 5.53035e-315
0
10 Buffer 3S~
219 2209 271 0 3 22
0 90 72 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U58D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 37 0
1 U
6748 0 0
2
5.89615e-315 5.531e-315
0
10 Buffer 3S~
219 2329 268 0 3 22
0 89 71 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U59A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 38 0
1 U
7393 0 0
2
5.89615e-315 5.53164e-315
0
10 Buffer 3S~
219 2441 269 0 3 22
0 88 69 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U59B
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 38 0
1 U
7699 0 0
2
5.89615e-315 5.53229e-315
0
10 Buffer 3S~
219 2563 266 0 3 22
0 87 68 86
0
0 0 112 270
8 BUFFER3S
-27 -51 29 -43
4 U59C
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 38 0
1 U
6638 0 0
2
5.89615e-315 5.53294e-315
0
10 Buffer 3S~
219 1695 666 0 3 22
0 86 58 66
0
0 0 112 512
8 BUFFER3S
-27 -51 29 -43
4 U59D
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 38 0
1 U
4595 0 0
2
5.89615e-315 5.53359e-315
0
9 2-In AND~
219 1909 878 0 3 22
0 49 85 61
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U47D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
9395 0 0
2
5.89615e-315 5.53423e-315
0
9 2-In AND~
219 859 456 0 3 22
0 61 84 145
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U51A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
3303 0 0
2
5.89615e-315 5.53488e-315
0
9 2-In AND~
219 961 457 0 3 22
0 61 83 143
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U51B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
4498 0 0
2
5.89615e-315 5.53553e-315
0
9 2-In AND~
219 1069 452 0 3 22
0 61 81 142
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U51C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
9728 0 0
2
5.89615e-315 5.53618e-315
0
9 2-In AND~
219 1185 452 0 3 22
0 61 82 144
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U51D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
3789 0 0
2
5.89615e-315 5.53682e-315
0
9 2-In AND~
219 1288 448 0 3 22
0 61 80 141
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U52A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
3978 0 0
2
5.89615e-315 5.53747e-315
0
9 2-In AND~
219 1504 446 0 3 22
0 61 79 139
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U52B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
3494 0 0
2
5.89615e-315 5.53812e-315
0
9 2-In AND~
219 1396 445 0 3 22
0 61 78 140
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U52C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
3507 0 0
2
5.89615e-315 5.53877e-315
0
9 2-In AND~
219 1612 446 0 3 22
0 61 77 115
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U52D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 31 0
1 U
5151 0 0
2
5.89615e-315 5.53941e-315
0
9 2-In AND~
219 1715 454 0 3 22
0 61 76 138
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U53A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
3701 0 0
2
5.89615e-315 5.54006e-315
0
9 2-In AND~
219 1826 447 0 3 22
0 61 75 137
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U53B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
8585 0 0
2
5.89615e-315 5.54071e-315
0
9 2-In AND~
219 1932 444 0 3 22
0 61 74 136
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U53C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
8809 0 0
2
5.89615e-315 5.54136e-315
0
9 2-In AND~
219 2041 440 0 3 22
0 61 73 135
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U53D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
5993 0 0
2
5.89615e-315 5.542e-315
0
9 2-In AND~
219 2154 446 0 3 22
0 61 72 134
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U54A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
8654 0 0
2
5.89615e-315 5.54265e-315
0
9 2-In AND~
219 2274 441 0 3 22
0 61 71 133
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U54B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
7223 0 0
2
5.89615e-315 5.5433e-315
0
9 2-In AND~
219 2386 447 0 3 22
0 61 69 132
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U54C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 33 0
1 U
3641 0 0
2
5.89615e-315 5.54395e-315
0
9 2-In AND~
219 2508 434 0 3 22
0 61 68 131
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U54D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 33 0
1 U
3104 0 0
2
5.89615e-315 5.54459e-315
0
10 Buffer 3S~
219 2051 266 0 3 22
0 67 135 13
0
0 0 112 602
8 BUFFER3S
-27 -51 29 -43
4 U55A
-13 -61 15 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
3296 0 0
2
5.89615e-315 5.54524e-315
0
10 TURING CPU
94 1181 745 0 17 35
0 57 56 55 2 48 47 51 54 53
52 55 56 66 57 50 49 4
10 TURING CPU
2 0 4240 0
0
3 U60
-14 -94 7 -86
0
0
0
0
0
0
35

0 6 7 8 9 10 11 12 13 14
15 26 27 28 29 37 38 0 6 7
8 9 10 11 12 13 14 15 26 27
28 29 37 38 0 0
0 0 0 0 1 0 0 0
1 U
8534 0 0
2
41410.4 44
0
5 CLOCK
94 494 660 0 3 5
0 49 50 42
5 CLOCK
3 0 4240 0
0
3 U62
-12 -44 9 -36
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
949 0 0
2
41410.4 45
0
4 BUSY
94 913 727 0 11 23
0 2 54 53 52 51 47 48 2 55
56 57
4 BUSY
4 0 4240 0
0
3 U61
-11 -56 10 -48
0
0
0
0
0
0
23

0 1 2 3 4 5 7 8 9 10
11 12 1 2 3 4 5 7 8 9
10 11 12 0
0 0 0 0 1 0 0 0
1 U
3371 0 0
2
5.8961e-315 0
0
398
0 0 3 0 0 4224 0 0 0 0 0 2
586 1190
609 1190
2 17 4 0 0 4224 0 22 194 0 0 3
1095 860
1140 860
1140 829
3 0 5 0 0 8320 0 42 0 0 300 4
305 437
305 1037
2759 1037
2759 741
3 0 6 0 0 8320 0 41 0 0 303 4
326 437
326 1039
2706 1039
2706 733
3 0 7 0 0 8320 0 40 0 0 213 4
347 437
347 1041
2652 1041
2652 729
0 3 8 0 0 8320 0 0 43 297 0 4
2810 745
2810 1035
284 1035
284 437
3 3 9 0 0 8320 0 39 108 0 0 4
638 151
638 276
2517 276
2517 247
3 3 10 0 0 8320 0 38 107 0 0 4
614 151
614 275
2396 275
2396 248
3 3 11 0 0 8320 0 37 106 0 0 4
591 151
591 276
2284 276
2284 246
3 3 12 0 0 8320 0 36 105 0 0 4
566 151
566 276
2164 276
2164 248
3 3 13 0 0 8320 0 35 193 0 0 4
543 151
543 275
2051 275
2051 251
3 3 14 0 0 8320 0 34 104 0 0 4
520 150
520 275
1942 275
1942 249
3 3 15 0 0 8320 0 33 103 0 0 4
499 150
499 275
1836 275
1836 246
3 3 16 0 0 8320 0 32 102 0 0 4
477 151
477 275
1726 275
1726 250
3 3 17 0 0 8320 0 31 101 0 0 4
453 151
453 275
1623 275
1623 246
3 3 18 0 0 8320 0 30 100 0 0 4
431 151
431 275
1515 275
1515 246
3 3 19 0 0 8320 0 29 99 0 0 4
409 150
409 276
1406 276
1406 245
3 3 20 0 0 8320 0 28 98 0 0 4
386 150
386 276
1298 276
1298 247
3 3 21 0 0 8320 0 27 97 0 0 4
364 150
364 276
1194 276
1194 247
3 3 22 0 0 8320 0 26 96 0 0 4
340 151
340 276
1079 276
1079 247
3 3 23 0 0 8320 0 25 95 0 0 4
316 152
316 275
974 275
974 247
3 3 24 0 0 8320 0 24 94 0 0 4
292 152
292 276
871 276
871 252
0 2 25 0 0 8192 0 0 43 56 0 3
272 421
272 422
295 422
2 2 25 0 0 4096 0 38 39 0 0 2
625 136
649 136
2 2 25 0 0 0 0 37 38 0 0 2
602 136
625 136
2 2 25 0 0 4096 0 36 37 0 0 2
577 136
602 136
2 2 25 0 0 0 0 35 36 0 0 2
554 136
577 136
2 2 25 0 0 0 0 34 35 0 0 4
531 135
544 135
544 136
554 136
2 2 25 0 0 0 0 33 34 0 0 2
510 135
531 135
2 2 25 0 0 0 0 32 33 0 0 3
488 136
488 135
510 135
2 2 25 0 0 0 0 31 32 0 0 2
464 136
488 136
2 2 25 0 0 0 0 30 31 0 0 2
442 136
464 136
2 2 25 0 0 0 0 29 30 0 0 3
420 135
420 136
442 136
2 2 25 0 0 0 0 28 29 0 0 4
397 135
397 136
420 136
420 135
2 2 25 0 0 0 0 27 28 0 0 4
375 135
375 136
397 136
397 135
2 2 25 0 0 0 0 26 27 0 0 3
351 136
375 136
375 135
2 2 25 0 0 0 0 25 26 0 0 3
327 137
327 136
351 136
2 2 25 0 0 0 0 24 25 0 0 2
303 137
327 137
1 1 26 0 0 4224 0 39 15 0 0 2
638 121
638 123
1 1 27 0 0 4224 0 38 14 0 0 2
614 121
614 123
1 1 28 0 0 4224 0 37 13 0 0 4
591 121
591 120
591 120
591 121
1 1 29 0 0 4224 0 36 12 0 0 2
566 121
566 122
1 1 30 0 0 4224 0 35 11 0 0 4
543 121
543 120
543 120
543 121
1 1 31 0 0 4224 0 34 10 0 0 2
520 120
520 123
1 1 32 0 0 4224 0 33 9 0 0 4
499 120
499 122
498 122
498 123
1 1 33 0 0 4224 0 32 8 0 0 3
477 121
477 124
476 124
1 1 34 0 0 4224 0 31 7 0 0 2
453 121
453 124
1 1 35 0 0 4224 0 30 6 0 0 2
431 121
431 124
1 1 36 0 0 8320 0 29 16 0 0 3
409 120
410 120
410 125
1 1 37 0 0 4224 0 28 5 0 0 2
386 120
386 124
1 1 38 0 0 4224 0 27 4 0 0 3
364 120
364 123
363 123
1 1 39 0 0 4224 0 26 3 0 0 2
340 121
340 125
1 1 40 0 0 4224 0 25 2 0 0 2
316 122
316 126
1 1 41 0 0 4224 0 24 1 0 0 2
292 122
292 126
1 0 42 0 0 8192 0 23 0 0 64 3
271 583
272 583
272 662
2 2 25 0 0 8320 0 24 23 0 0 4
303 137
272 137
272 547
271 547
2 2 25 0 0 0 0 41 40 0 0 2
337 422
358 422
2 2 25 0 0 0 0 42 41 0 0 2
316 422
337 422
2 2 25 0 0 0 0 43 42 0 0 2
295 422
316 422
1 1 43 0 0 4224 0 40 17 0 0 4
347 407
347 408
348 408
348 409
1 1 44 0 0 4224 0 41 20 0 0 3
326 407
327 407
327 408
1 1 45 0 0 4224 0 42 19 0 0 2
305 407
305 410
1 1 46 0 0 4224 0 43 18 0 0 4
284 407
284 408
283 408
283 409
1 3 42 0 0 12288 0 21 195 0 0 4
246 664
272 664
272 662
455 662
6 6 47 0 0 4224 0 194 196 0 0 2
1098 754
946 754
7 5 48 0 0 4224 0 196 194 0 0 2
946 745
1098 745
4 8 2 0 0 4224 0 194 196 0 0 2
1098 736
946 736
1 16 49 0 0 4096 0 195 194 0 0 2
518 671
1199 671
2 15 50 0 0 20480 0 195 194 0 0 7
518 662
526 662
526 643
699 643
699 644
1208 644
1208 671
0 1 42 0 0 8320 0 0 22 64 0 3
436 662
436 860
1059 860
1 1 2 0 0 0 0 196 44 0 0 2
880 709
787 709
5 7 51 0 0 12416 0 196 194 0 0 4
880 745
842 745
842 799
1098 799
10 4 52 0 0 4224 0 194 196 0 0 4
1098 790
851 790
851 736
880 736
3 9 53 0 0 12416 0 196 194 0 0 4
880 727
857 727
857 781
1098 781
8 2 54 0 0 4224 0 194 196 0 0 4
1098 772
866 772
866 718
880 718
3 9 55 0 0 4096 0 194 196 0 0 2
1098 727
946 727
2 10 56 0 0 4096 0 194 196 0 0 2
1098 718
946 718
1 11 57 0 0 4096 0 194 196 0 0 2
1098 709
946 709
14 1 57 0 0 4224 0 194 136 0 0 4
1257 718
1595 718
1595 713
1680 713
12 1 56 0 0 4224 0 194 137 0 0 4
1257 728
1598 728
1598 771
1680 771
2 0 58 0 0 8320 0 158 0 0 86 3
2173 816
2173 841
1695 841
2 2 58 0 0 0 0 157 158 0 0 2
2173 766
2173 816
2 2 58 0 0 0 0 155 157 0 0 2
2173 712
2173 766
2 2 58 0 0 0 0 156 155 0 0 2
2173 660
2173 712
1 11 55 0 0 12416 0 138 194 0 0 4
1680 822
1592 822
1592 740
1257 740
3 2 58 0 0 0 0 139 138 0 0 2
1695 856
1695 833
0 3 59 0 0 8320 0 0 136 135 0 3
1743 701
1743 713
1710 713
2 2 60 0 0 4224 0 149 148 0 0 2
1761 665
1761 668
3 0 61 0 0 4224 0 176 0 0 111 2
1908 854
1908 483
2 2 62 0 0 4224 0 146 147 0 0 2
2285 823
2284 823
2 2 63 0 0 4224 0 145 142 0 0 2
2282 773
2281 773
2 2 64 0 0 4224 0 143 141 0 0 2
2280 718
2279 718
2 2 65 0 0 4224 0 144 140 0 0 2
2278 667
2277 667
0 0 50 0 0 0 0 0 0 223 69 4
886 960
886 961
699 961
699 644
1 13 66 0 0 12416 0 133 194 0 0 4
1641 666
1597 666
1597 707
1257 707
0 0 49 0 0 0 0 0 0 224 68 3
887 917
718 917
718 671
1 0 67 0 0 4096 0 193 0 0 331 2
2051 281
2051 297
0 3 13 0 0 0 0 0 193 99 0 2
2051 242
2051 251
1 1 13 0 0 0 0 79 81 0 0 3
2067 242
2049 242
2049 211
1 0 61 0 0 0 0 192 0 0 102 3
2498 455
2498 483
2376 483
2 5 68 0 0 8192 0 192 0 0 152 7
2516 455
2530 455
2530 408
2552 408
2552 406
2551 406
2551 403
1 0 61 0 0 0 0 191 0 0 105 3
2376 468
2376 483
2264 483
2 5 69 0 0 8192 0 191 116 0 0 7
2394 468
2408 468
2408 421
2430 421
2430 419
2429 419
2429 416
1 0 70 0 0 4096 0 116 0 0 295 2
2416 461
2416 534
1 0 61 0 0 0 0 190 0 0 107 3
2264 462
2264 483
2144 483
2 5 71 0 0 8192 0 190 0 0 156 7
2282 462
2296 462
2296 415
2318 415
2318 413
2317 413
2317 411
1 0 61 0 0 0 0 189 0 0 109 3
2144 467
2144 483
2031 483
2 5 72 0 0 8192 0 189 0 0 158 6
2162 467
2176 467
2176 420
2198 420
2198 418
2197 418
1 0 61 0 0 0 0 188 0 0 111 3
2031 461
2031 483
1922 483
2 5 73 0 0 8192 0 188 0 0 160 5
2049 461
2061 461
2061 415
2083 415
2083 414
1 0 61 0 0 0 0 187 0 0 113 3
1922 465
1922 483
1816 483
2 0 74 0 0 8192 0 187 0 0 162 4
1940 465
1952 465
1952 414
1976 414
1 0 61 0 0 0 0 186 0 0 115 3
1816 468
1816 483
1705 483
2 5 75 0 0 8192 0 186 0 0 164 4
1834 468
1846 468
1846 417
1869 417
1 0 61 0 0 0 0 185 0 0 117 3
1705 475
1705 483
1602 483
2 5 76 0 0 8192 0 185 0 0 166 4
1723 475
1738 475
1738 426
1761 426
1 0 61 0 0 0 0 184 0 0 121 3
1602 467
1602 483
1493 483
2 5 77 0 0 8192 0 184 0 0 168 4
1620 467
1635 467
1635 421
1658 421
1 0 61 0 0 0 0 183 0 0 123 3
1386 466
1386 483
1278 483
2 5 78 0 0 8192 0 183 0 0 172 4
1404 466
1417 466
1417 421
1440 421
1 0 61 0 0 0 0 182 0 0 119 5
1494 467
1494 475
1493 475
1493 483
1386 483
2 5 79 0 0 8192 0 182 0 0 170 4
1512 467
1527 467
1527 421
1550 421
1 0 61 0 0 0 0 181 0 0 126 3
1278 469
1278 483
1175 483
2 5 80 0 0 8192 0 181 0 0 176 4
1296 469
1309 469
1309 424
1332 424
2 5 81 0 0 8192 0 179 112 0 0 5
1077 473
1091 473
1091 429
1111 429
1111 428
1 0 61 0 0 0 0 180 0 0 0 3
1175 473
1175 483
839 483
2 5 82 0 0 8192 0 180 0 0 174 4
1193 473
1204 473
1204 428
1227 428
1 0 61 0 0 0 0 179 0 0 126 2
1059 473
1059 483
1 0 61 0 0 0 0 178 0 0 126 4
951 478
951 473
951 473
951 483
2 5 83 0 0 8192 0 178 111 0 0 5
969 478
981 478
981 433
1005 433
1005 432
0 1 61 0 0 0 0 0 177 126 0 2
849 483
849 477
2 0 84 0 0 8192 0 177 0 0 183 4
867 477
879 477
879 430
900 430
2 0 85 0 0 4096 0 176 0 0 222 2
1917 899
1917 967
1 0 49 0 0 0 0 176 0 0 224 2
1899 899
1899 908
1 1 59 0 0 0 0 149 148 0 0 3
1761 701
1743 701
1743 668
2 2 58 0 0 0 0 136 175 0 0 2
1695 724
1695 677
1 3 86 0 0 8192 0 175 161 0 0 6
1710 666
1710 619
832 619
832 334
1122 334
1122 286
3 0 86 0 0 0 0 163 0 0 150 2
1238 285
1238 334
3 0 86 0 0 0 0 162 0 0 150 2
1343 285
1343 334
3 0 86 0 0 0 0 164 0 0 150 2
1451 283
1451 334
3 0 86 0 0 0 0 165 0 0 150 2
1561 283
1561 334
3 0 86 0 0 0 0 166 0 0 150 2
1669 283
1669 334
3 0 86 0 0 0 0 167 0 0 150 2
1772 286
1772 334
3 0 86 0 0 0 0 168 0 0 150 2
1880 283
1880 334
3 0 86 0 0 0 0 169 0 0 150 2
1987 287
1987 334
3 0 86 0 0 0 0 170 0 0 150 2
2094 286
2094 334
3 0 86 0 0 0 0 171 0 0 150 2
2208 287
2208 334
3 0 86 0 0 0 0 172 0 0 150 2
2328 284
2328 334
3 0 86 0 0 0 0 173 0 0 150 2
2440 285
2440 334
0 3 86 0 0 4224 0 0 174 137 0 3
1122 334
2562 334
2562 282
4 1 87 0 0 41088 0 0 174 363 0 11
2517 160
2518 160
2518 159
2517 159
2517 161
2516 161
2516 161
2529 161
2529 144
2562 144
2562 252
2 5 68 0 0 4224 0 174 123 0 0 2
2551 267
2551 406
4 1 88 0 0 36992 0 0 173 359 0 10
2396 163
2396 162
2395 162
2395 164
2394 164
2394 162
2407 162
2407 147
2440 147
2440 255
2 5 69 0 0 4224 0 173 116 0 0 2
2429 270
2429 416
4 1 89 0 0 36992 0 0 172 355 0 10
2284 162
2284 161
2283 161
2283 163
2282 163
2282 162
2295 162
2295 146
2328 146
2328 254
2 5 71 0 0 4224 0 172 124 0 0 2
2317 269
2317 411
4 1 90 0 0 28800 0 0 171 351 0 8
2163 164
2163 166
2162 166
2162 166
2175 166
2175 149
2208 149
2208 257
2 5 72 0 0 4224 0 171 120 0 0 2
2197 272
2197 418
4 1 91 0 0 28800 0 0 170 347 0 8
2049 163
2049 165
2048 165
2048 162
2061 162
2061 148
2094 148
2094 256
2 5 73 0 0 4224 0 170 118 0 0 2
2083 271
2083 414
4 1 92 0 0 28800 0 0 169 345 0 8
1942 165
1942 166
1941 166
1941 165
1954 165
1954 149
1987 149
1987 257
2 5 74 0 0 4224 0 169 117 0 0 2
1976 272
1976 416
4 1 93 0 0 24704 0 0 168 367 0 7
1836 162
1834 162
1834 161
1847 161
1847 145
1880 145
1880 253
2 5 75 0 0 4224 0 168 119 0 0 2
1869 268
1869 418
4 1 94 0 0 20608 0 0 167 394 0 6
1726 163
1726 162
1739 162
1739 148
1772 148
1772 256
2 5 76 0 0 4224 0 167 122 0 0 2
1761 271
1761 426
4 1 95 0 0 20608 0 0 166 398 0 6
1623 163
1623 164
1636 164
1636 145
1669 145
1669 253
2 5 77 0 0 4224 0 166 121 0 0 2
1658 268
1658 421
4 1 96 0 0 20608 0 0 165 390 0 6
1515 163
1515 164
1528 164
1528 145
1561 145
1561 253
2 5 79 0 0 4224 0 165 115 0 0 2
1550 268
1550 423
4 1 97 0 0 16512 0 0 164 386 0 5
1406 163
1418 163
1418 145
1451 145
1451 253
2 5 78 0 0 4224 0 164 113 0 0 2
1440 268
1440 426
4 1 98 0 0 16512 0 0 163 379 0 5
1194 164
1205 164
1205 147
1238 147
1238 255
2 5 82 0 0 4224 0 163 110 0 0 2
1227 270
1227 428
4 1 99 0 0 16512 0 0 162 383 0 5
1298 163
1310 163
1310 147
1343 147
1343 255
2 5 80 0 0 4224 0 162 114 0 0 2
1332 270
1332 426
4 1 100 0 0 20608 0 54 161 0 0 6
1079 165
1079 166
1089 166
1089 148
1122 148
1122 256
3 0 86 0 0 0 0 160 0 0 137 2
1016 284
1016 334
3 0 86 0 0 0 0 159 0 0 137 2
911 285
911 334
1 3 66 0 0 0 0 133 175 0 0 2
1641 666
1680 666
2 5 81 0 0 4224 0 161 112 0 0 2
1111 271
1111 428
2 5 83 0 0 4224 0 160 111 0 0 2
1005 269
1005 432
2 5 84 0 0 4224 0 159 109 0 0 2
900 270
900 433
4 1 101 0 0 16512 0 48 160 0 0 5
974 164
983 164
983 149
1016 149
1016 254
4 1 102 0 0 16512 0 51 159 0 0 5
871 167
882 167
882 152
911 152
911 255
1 0 103 0 0 4096 0 144 0 0 189 2
2242 667
2242 649
3 1 104 0 0 4224 0 158 147 0 0 2
2188 805
2284 805
3 1 105 0 0 4224 0 157 142 0 0 2
2188 755
2281 755
3 1 103 0 0 4224 0 156 140 0 0 2
2188 649
2277 649
3 1 106 0 0 4224 0 155 141 0 0 4
2188 701
2244 701
2244 700
2279 700
10 1 107 0 0 8320 0 45 156 0 0 4
2077 737
2125 737
2125 649
2158 649
1 0 104 0 0 0 0 146 0 0 187 3
2249 823
2248 823
2248 805
7 1 108 0 0 4224 0 45 158 0 0 4
2077 765
2127 765
2127 805
2158 805
4 1 109 0 0 4224 0 147 153 0 0 2
2332 805
2358 805
1 0 105 0 0 0 0 145 0 0 188 3
2246 773
2245 773
2245 755
1 0 106 0 0 0 0 143 0 0 190 2
2244 718
2244 700
9 1 110 0 0 4224 0 45 155 0 0 4
2077 747
2129 747
2129 701
2158 701
4 0 111 0 0 12288 0 45 0 0 290 5
1981 753
1970 753
1970 597
2601 597
2601 501
3 0 112 0 0 12288 0 45 0 0 292 5
1981 744
1973 744
1973 600
2607 600
2607 513
2 0 113 0 0 12288 0 45 0 0 294 5
1981 735
1977 735
1977 603
2612 603
2612 526
1 0 114 0 0 12288 0 45 0 0 296 5
1981 727
1980 727
1980 606
2617 606
2617 541
2 3 115 0 0 4224 0 101 184 0 0 4
1612 261
1612 400
1611 400
1611 422
2 0 116 0 0 4096 0 154 0 0 225 2
2382 904
2382 932
1 0 50 0 0 0 0 154 0 0 223 2
2364 904
2364 946
2 3 117 0 0 4096 0 153 154 0 0 2
2373 816
2373 859
2 2 117 0 0 0 0 152 153 0 0 4
2371 766
2371 801
2373 801
2373 816
2 2 117 0 0 4224 0 151 152 0 0 2
2371 711
2371 766
2 2 117 0 0 0 0 150 151 0 0 2
2371 660
2371 711
4 1 118 0 0 4224 0 142 152 0 0 2
2329 755
2356 755
4 1 119 0 0 4224 0 141 151 0 0 2
2327 700
2356 700
4 1 120 0 0 4224 0 140 150 0 0 2
2325 649
2356 649
1 0 7 0 0 0 0 126 0 0 213 2
2670 620
2652 620
1 3 7 0 0 0 0 125 150 0 0 5
2652 589
2652 732
2406 732
2406 649
2386 649
8 1 121 0 0 4224 0 45 157 0 0 2
2077 755
2158 755
0 4 67 0 0 12288 0 0 148 331 0 5
871 298
827 298
827 612
1743 612
1743 620
3 5 122 0 0 4224 0 137 45 0 0 2
1710 771
1981 771
2 0 85 0 0 0 0 139 0 0 222 2
1704 901
1704 967
1 0 116 0 0 4096 0 139 0 0 225 2
1686 901
1686 932
2 2 58 0 0 0 0 137 138 0 0 2
1695 782
1695 833
2 2 58 0 0 0 0 136 137 0 0 2
1695 724
1695 782
3 6 123 0 0 8320 0 138 45 0 0 3
1710 822
1710 779
1981 779
2 0 85 0 0 4224 0 134 0 0 0 2
937 967
2395 967
1 0 50 0 0 12416 0 134 0 0 0 4
901 967
886 967
886 946
2394 946
1 0 49 0 0 12416 0 135 0 0 0 4
896 932
887 932
887 908
2394 908
2 0 116 0 0 4224 0 135 0 0 0 2
932 932
2393 932
4 0 111 0 0 0 0 123 0 0 290 4
2565 451
2565 486
2566 486
2566 501
4 0 111 0 0 0 0 116 0 0 290 2
2443 461
2443 501
4 0 111 0 0 0 0 124 0 0 290 2
2331 456
2331 501
4 0 111 0 0 0 0 120 0 0 290 2
2211 463
2211 501
4 0 111 0 0 0 0 118 0 0 290 2
2097 459
2097 501
4 0 111 0 0 0 0 117 0 0 290 4
1990 461
1990 486
1989 486
1989 501
4 0 111 0 0 0 0 119 0 0 290 2
1883 463
1883 501
4 0 111 0 0 0 0 122 0 0 290 2
1775 471
1775 501
4 0 124 0 0 12288 0 121 0 0 289 4
1672 466
1672 479
1671 479
1671 493
4 0 124 0 0 4096 0 115 0 0 289 2
1564 468
1564 493
4 0 124 0 0 0 0 113 0 0 289 4
1454 471
1454 479
1453 479
1453 493
4 0 124 0 0 0 0 114 0 0 289 4
1346 471
1346 481
1345 481
1345 493
4 0 124 0 0 0 0 110 0 0 289 2
1241 473
1241 493
4 0 124 0 0 0 0 112 0 0 289 2
1125 473
1125 493
4 0 124 0 0 0 0 111 0 0 289 2
1019 477
1019 493
3 0 112 0 0 0 0 123 0 0 292 4
2556 451
2556 498
2555 498
2555 513
3 0 112 0 0 0 0 116 0 0 292 4
2434 461
2434 498
2433 498
2433 513
3 0 112 0 0 0 0 124 0 0 292 2
2322 456
2322 513
3 0 112 0 0 0 0 120 0 0 292 4
2202 463
2202 498
2201 498
2201 513
3 0 125 0 0 4096 0 118 0 0 291 2
2088 459
2088 507
3 0 125 0 0 0 0 117 0 0 291 2
1981 461
1981 507
3 0 125 0 0 0 0 119 0 0 291 4
1874 463
1874 492
1873 492
1873 507
3 0 125 0 0 0 0 122 0 0 291 2
1766 471
1766 507
3 0 112 0 0 0 0 121 0 0 292 2
1663 466
1663 513
3 0 112 0 0 0 0 115 0 0 292 2
1555 468
1555 513
3 0 112 0 0 0 0 113 0 0 292 2
1445 471
1445 513
3 0 112 0 0 0 0 114 0 0 292 2
1337 471
1337 513
3 0 125 0 0 0 0 110 0 0 291 2
1232 473
1232 507
3 0 125 0 0 0 0 112 0 0 291 4
1116 473
1116 492
1115 492
1115 507
3 0 125 0 0 0 0 111 0 0 291 2
1010 477
1010 507
2 0 113 0 0 0 0 123 0 0 294 2
2547 451
2547 526
2 0 113 0 0 0 0 116 0 0 294 2
2425 461
2425 526
2 0 126 0 0 4096 0 124 0 0 293 2
2313 456
2313 519
2 0 126 0 0 0 0 120 0 0 293 2
2193 463
2193 519
2 0 113 0 0 0 0 118 0 0 294 4
2079 459
2079 511
2078 511
2078 526
2 0 113 0 0 0 0 117 0 0 294 2
1972 461
1972 526
2 0 126 0 0 0 0 119 0 0 293 2
1865 463
1865 519
2 0 126 0 0 0 0 122 0 0 293 2
1757 471
1757 519
2 0 113 0 0 0 0 121 0 0 294 2
1654 466
1654 526
2 0 113 0 0 0 0 115 0 0 294 2
1546 468
1546 526
2 0 126 0 0 0 0 113 0 0 293 2
1436 471
1436 519
2 0 126 0 0 0 0 114 0 0 293 2
1328 471
1328 519
2 0 113 0 0 0 0 110 0 0 294 2
1223 473
1223 526
2 0 113 0 0 0 0 112 0 0 294 2
1107 473
1107 526
2 0 126 0 0 0 0 111 0 0 293 2
1001 477
1001 519
1 0 114 0 0 0 0 123 0 0 296 2
2538 451
2538 541
1 0 114 0 0 0 0 124 0 0 296 4
2304 456
2304 526
2303 526
2303 541
1 0 70 0 0 0 0 120 0 0 295 2
2184 463
2184 534
1 0 114 0 0 0 0 118 0 0 296 2
2070 459
2070 541
1 0 70 0 0 0 0 117 0 0 295 2
1963 461
1963 534
1 0 114 0 0 0 0 119 0 0 296 2
1856 463
1856 541
1 0 70 0 0 0 0 122 0 0 295 2
1748 471
1748 534
1 0 114 0 0 0 0 121 0 0 296 2
1645 466
1645 541
1 0 70 0 0 0 0 115 0 0 295 2
1537 468
1537 534
1 0 114 0 0 0 0 113 0 0 296 2
1427 471
1427 541
1 0 70 0 0 0 0 114 0 0 295 2
1319 471
1319 534
1 0 114 0 0 0 0 110 0 0 296 2
1214 473
1214 541
1 0 70 0 0 0 0 112 0 0 295 4
1098 473
1098 519
1097 519
1097 534
1 0 114 0 0 0 0 111 0 0 296 2
992 477
992 541
4 0 124 0 0 0 0 109 0 0 289 2
914 478
914 493
3 0 125 0 0 0 0 109 0 0 291 2
905 478
905 507
2 0 126 0 0 0 0 109 0 0 293 2
896 478
896 519
1 0 70 0 0 0 0 109 0 0 295 2
887 478
887 534
3 0 124 0 0 8320 0 132 0 0 0 3
2828 532
2828 493
839 493
4 0 111 0 0 8320 0 132 0 0 0 3
2810 538
2810 501
838 501
3 0 125 0 0 8320 0 129 0 0 0 3
2777 533
2777 507
838 507
4 0 112 0 0 8320 0 129 0 0 0 3
2759 539
2759 513
838 513
3 0 126 0 0 8320 0 128 0 0 0 3
2724 533
2724 519
839 519
4 0 113 0 0 8320 0 128 0 0 0 3
2706 539
2706 526
839 526
3 0 70 0 0 8320 0 125 0 0 0 3
2670 535
2670 534
839 534
4 0 114 0 0 4224 0 125 0 0 0 2
2652 541
840 541
0 3 8 0 0 0 0 0 153 298 0 5
2810 617
2810 746
2407 746
2407 805
2388 805
1 1 8 0 0 0 0 132 131 0 0 3
2810 586
2810 617
2828 617
2 2 127 0 0 4224 0 131 132 0 0 2
2828 581
2828 586
0 3 5 0 0 0 0 0 152 301 0 5
2759 618
2759 741
2405 741
2405 755
2386 755
1 1 5 0 0 0 0 129 130 0 0 3
2759 587
2759 618
2777 618
2 2 128 0 0 4224 0 130 129 0 0 2
2777 582
2777 587
0 3 6 0 0 0 0 0 151 304 0 5
2706 618
2706 736
2403 736
2403 700
2386 700
1 1 6 0 0 0 0 128 127 0 0 3
2706 587
2706 618
2724 618
2 2 129 0 0 4224 0 127 128 0 0 2
2724 582
2724 587
2 2 130 0 0 4224 0 126 125 0 0 2
2670 584
2670 589
2 3 131 0 0 4224 0 108 192 0 0 4
2506 262
2506 347
2507 347
2507 410
2 3 132 0 0 20608 0 107 191 0 0 6
2385 263
2385 278
2386 278
2386 347
2385 347
2385 423
2 3 133 0 0 4224 0 106 190 0 0 2
2273 261
2273 417
2 3 134 0 0 4224 0 105 189 0 0 2
2153 263
2153 422
2 3 135 0 0 4224 0 193 188 0 0 2
2040 266
2040 416
2 3 136 0 0 4224 0 104 187 0 0 2
1931 264
1931 420
2 3 137 0 0 4224 0 103 186 0 0 2
1825 261
1825 423
2 3 138 0 0 12416 0 102 185 0 0 4
1715 265
1715 339
1714 339
1714 430
2 3 139 0 0 12416 0 100 182 0 0 4
1504 261
1504 340
1503 340
1503 422
2 3 140 0 0 4224 0 99 183 0 0 2
1395 260
1395 421
2 3 141 0 0 4224 0 98 181 0 0 2
1287 262
1287 424
2 3 142 0 0 4224 0 96 179 0 0 2
1068 262
1068 428
2 3 143 0 0 8320 0 95 178 0 0 3
963 262
960 262
960 433
2 3 144 0 0 12416 0 97 180 0 0 4
1183 262
1183 343
1184 343
1184 428
2 3 145 0 0 8320 0 94 177 0 0 3
860 267
858 267
858 432
2 0 136 0 0 0 0 104 0 0 0 4
1931 264
1931 265
1931 265
1931 264
3 0 19 0 0 0 0 99 0 0 384 2
1406 245
1406 241
3 0 21 0 0 0 0 97 0 0 377 2
1194 247
1194 242
3 0 22 0 0 0 0 96 0 0 374 2
1079 247
1079 241
3 0 23 0 0 0 0 95 0 0 368 2
974 247
974 241
0 3 24 0 0 0 0 0 94 371 0 2
871 246
871 252
1 0 67 0 0 0 0 108 0 0 331 3
2517 277
2517 297
2164 297
1 0 67 0 0 0 0 107 0 0 328 2
2396 278
2396 297
1 0 67 0 0 0 0 106 0 0 328 2
2284 276
2284 297
1 1 67 0 0 8320 0 105 94 0 0 6
2164 278
2164 297
1199 297
1199 298
871 298
871 282
1 0 67 0 0 0 0 104 0 0 331 2
1942 279
1942 297
1 0 67 0 0 0 0 103 0 0 331 2
1836 276
1836 297
1 0 67 0 0 0 0 102 0 0 331 2
1726 280
1726 297
1 0 67 0 0 0 0 101 0 0 331 2
1623 276
1623 297
1 0 67 0 0 0 0 100 0 0 331 2
1515 276
1515 297
1 0 67 0 0 0 0 99 0 0 331 2
1406 275
1406 297
1 0 67 0 0 0 0 98 0 0 331 2
1298 277
1298 297
1 0 67 0 0 0 0 97 0 0 331 2
1194 277
1194 297
1 0 67 0 0 0 0 96 0 0 331 2
1079 277
1079 297
1 0 67 0 0 0 0 95 0 0 331 2
974 277
974 297
0 3 14 0 0 0 0 0 104 343 0 2
1942 243
1942 249
1 1 14 0 0 0 0 76 78 0 0 3
1942 212
1942 243
1960 243
2 2 146 0 0 4224 0 78 76 0 0 2
1960 207
1960 212
1 4 92 0 0 0 0 77 76 0 0 2
1942 166
1942 164
2 2 147 0 0 4224 0 79 81 0 0 2
2067 206
2067 211
1 4 91 0 0 0 0 80 81 0 0 2
2049 165
2049 163
0 3 12 0 0 0 0 0 105 349 0 4
2163 243
2163 245
2164 245
2164 248
1 1 12 0 0 0 0 82 84 0 0 3
2163 212
2163 243
2181 243
2 2 148 0 0 4224 0 84 82 0 0 2
2181 207
2181 212
1 4 90 0 0 0 0 83 82 0 0 2
2163 166
2163 164
0 3 11 0 0 0 0 0 106 353 0 2
2284 241
2284 246
1 1 11 0 0 0 0 87 85 0 0 3
2284 210
2284 241
2302 241
2 2 149 0 0 4224 0 85 87 0 0 2
2302 205
2302 210
1 4 89 0 0 0 0 86 87 0 0 2
2284 164
2284 162
0 3 10 0 0 0 0 0 107 357 0 2
2396 241
2396 248
1 1 10 0 0 0 0 88 90 0 0 3
2396 210
2396 241
2414 241
2 2 150 0 0 4224 0 90 88 0 0 2
2414 205
2414 210
1 4 88 0 0 0 0 89 88 0 0 2
2396 164
2396 162
0 3 9 0 0 0 0 0 108 361 0 2
2517 239
2517 247
1 1 9 0 0 0 0 91 93 0 0 3
2517 208
2517 239
2535 239
2 2 151 0 0 4224 0 93 91 0 0 2
2535 203
2535 208
1 4 87 0 0 0 0 92 91 0 0 2
2517 162
2517 160
0 3 15 0 0 0 0 0 103 365 0 2
1836 240
1836 246
1 1 15 0 0 0 0 75 73 0 0 3
1836 209
1836 240
1854 240
2 2 152 0 0 4224 0 73 75 0 0 2
1854 204
1854 209
1 4 93 0 0 0 0 74 75 0 0 2
1836 163
1836 161
1 1 23 0 0 0 0 48 46 0 0 3
974 212
974 243
992 243
2 2 153 0 0 4224 0 46 48 0 0 2
992 207
992 212
1 4 101 0 0 0 0 47 48 0 0 2
974 166
974 164
1 1 24 0 0 0 0 51 49 0 0 3
871 215
871 246
889 246
2 2 154 0 0 4224 0 49 51 0 0 2
889 210
889 215
1 4 102 0 0 0 0 50 51 0 0 2
871 169
871 167
1 1 22 0 0 0 0 54 52 0 0 3
1079 213
1079 244
1097 244
2 2 155 0 0 4224 0 52 54 0 0 2
1097 208
1097 213
1 4 100 0 0 0 0 53 54 0 0 2
1079 167
1079 165
1 1 21 0 0 0 0 55 57 0 0 3
1194 212
1194 243
1212 243
2 2 156 0 0 4224 0 57 55 0 0 2
1212 207
1212 212
1 4 98 0 0 0 0 56 55 0 0 2
1194 166
1194 164
0 3 20 0 0 0 0 0 98 381 0 2
1298 241
1298 247
1 1 20 0 0 0 0 60 58 0 0 3
1298 210
1298 241
1316 241
2 2 157 0 0 4224 0 58 60 0 0 2
1316 205
1316 210
1 4 99 0 0 0 0 59 60 0 0 2
1298 164
1298 162
1 1 19 0 0 0 0 61 63 0 0 3
1406 210
1406 241
1424 241
2 2 158 0 0 4224 0 63 61 0 0 2
1424 205
1424 210
1 4 97 0 0 0 0 62 61 0 0 2
1406 164
1406 162
0 3 18 0 0 0 0 0 100 388 0 2
1515 241
1515 246
1 1 18 0 0 0 0 66 64 0 0 3
1515 210
1515 241
1533 241
2 2 159 0 0 4224 0 64 66 0 0 2
1533 205
1533 210
1 4 96 0 0 0 0 65 66 0 0 2
1515 164
1515 162
0 3 16 0 0 0 0 0 102 392 0 2
1726 242
1726 250
1 1 16 0 0 0 0 70 72 0 0 3
1726 211
1726 242
1744 242
2 2 160 0 0 4224 0 72 70 0 0 2
1744 206
1744 211
1 4 94 0 0 0 0 71 70 0 0 2
1726 165
1726 163
0 3 17 0 0 0 0 0 101 396 0 2
1623 242
1623 246
1 1 17 0 0 0 0 67 69 0 0 3
1623 211
1623 242
1641 242
2 2 161 0 0 4224 0 69 67 0 0 2
1641 206
1641 211
1 4 95 0 0 0 0 68 67 0 0 2
1623 165
1623 163
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 46
87 94 276 138
97 102 265 134
46 Configuraci�n inicial 
         de la cinta:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 44
79 368 260 412
89 376 249 408
44     Posici�n inicial 
        del cabezal:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
101 646 202 670
111 654 191 670
10 Start/Stop
-27 0 0 0 400 0 0 0 0 3 2 1 34
12 Arial Narrow
0 0 0 14
281 12 426 55
291 20 415 51
14 Inicializaci�n
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
2514 262 2751 286
2524 270 2740 286
27 << Este cable contiene a OB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
2516 282 2705 306
2526 290 2694 306
21 << Este contiene a IB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 166
2570 403 3031 467
2580 411 3020 459
166 <<De todos estos AND, solo el correspondiente a la pos 
actual estar� en 1, con lo que el FF correspondiente se 
conectara a los cables de entrada IB y  salida OB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 59
2691 612 3042 656
2711 628 3021 660
59 <<Este registro de 4B  almacena 
la pos actual del cabezal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
2566 129 2643 153
2576 137 2632 153
7 <<-Tape
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1700 874 1778 889
1714 885 1763 896
7 Step 00
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
2386 871 2464 886
2400 882 2449 893
7 Step 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1912 869 1992 884
1927 881 1976 892
7 Step 01
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
